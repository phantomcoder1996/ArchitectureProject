Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
Entity ROM is

port(
address: in std_logic_vector(6 downto 0);
dataout: out std_logic_vector(28 downto 0)

);

end entity;


Architecture ROMArch of ROM is

type romtype is Array(0 to 97) of std_logic_vector(28 downto 0);

signal rom:romtype:=
(
"00000100000000000000100000000",
"10001000000000000000000000000",
"00000000000001010001000000100",
"00000000000000000000000000000",
"00000110000101001000000011000",
"10000001001010000010100110000",
"00011001001000010010001110000",
"00000110000101000000000101000",
"10000000000100001000000010000",
"01011001001000000001001110000",
"00000000000000000000000000000",
"00000000000001110000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000011001100100100000101001",
"10000010001010100000000101010",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000110000100100000000101000",
"10000000011000001100000010010",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000110011100101100000011000",
"10000000000000000000000000010",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000111000100100000011100000",
"10001000000000000000000000010",
"00000000000000000000000000000",
"00000000000000000000000000000",
"01000001001000000101000110001",
"00000000000000000000000000000",
"00000000000000000000000000000",
"01000001001000001101001110000",
"00000110100100100010000101000",
"00000000001000001110001010000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000110100100101110000011000",
"00000000000000000010001000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"11100001001010000011000000000",
"00000000000000000010001000000",
"00000111100100100000011100000",
"10000010001010100010000101000",
"00000000000000000010001000000",
"00000011101000100100011100000",
"00000110000100100000000101000",
"10000000101000001100000010000",
"00000110000101100010000101000",
"00000000000000000010001000000",
"00000011101000100100011100000",
"00000110011100101100000011000",
"10000110000101100010000101000",
"00000000000000000010001000000",
"00000010001000101100001101000",
"00000011000100100000000101000",
"00100010100000100000001000000",
"00000011000100100000000101000",
"00100000011000001100001000000",
"00011011001000010000101100000",
"00100010101000101100001000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000110100100100000000101000",
"10000000001000001100000010011",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000110101100101100000011000",
"10000000000000000000000000011",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000000000000000000000000000",
"00000100000000000000100000000",
"10001000000000000000000000000",
"00000101100100100001010100000",
"10000000000000000000000000011",
"11100011001011100011000000000",
"00000000000000000010001000000",
"01100011000001100001001000000",
"00000111100100100001010100000",
"10000010001011100010000101000",
"00000000000000000010001000000"
);
begin

dataout<=rom(to_integer(unsigned(address)));

End ROMArch;
